Agent policy,Adversary policy,touches
maddpg,maddpg,1.014985014985015
maddpg,ddpg,1.1458541458541458
ddpg,maddpg,0.7542457542457542
ddpg,ddpg,0.6963036963036963
